module lab3();

endmodule;