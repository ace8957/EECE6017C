module mem(mclock, pclock, resetn, run, done, bus);
	
	input mclock, pclock, resetn, run;
	output done;
	output [8:0] bus;
	
	
	
endmodule